--romForwardZetas
--Used as ROM to store the forward NTT twiddle factors

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use IEEE.math_real.all;
use work.GlobalVars.all;

entity romForwardZetas is
  generic (
    width   : integer := 32;
    depth   : integer := 8
  );

  	PORT
	(
		address 		: IN STD_LOGIC_VECTOR (depth - 1 DOWNTO 0);
		clk		    : IN STD_LOGIC;
		q		        : OUT STD_LOGIC_VECTOR (width - 1 DOWNTO 0)
	);

  attribute RAM_STYLE         : string;
  attribute RAM_STYLE of romForwardZetas : entity is "block";
end entity;

architecture RTL of romForwardZetas is
  subtype word_t is std_logic_vector(width - 1 downto 0);
  type memory_t is array(0 to 2**depth - 1) of word_t;

  signal ram : memory_t := (
    0 => x"00000000",
    1 => x"000064F7",
    2 => x"00581103",
    3 => x"0077F504",
    4 => x"00039E44",
    5 => x"00740119",
    6 => x"00728129",
    7 => x"00071E24",
    8 => x"001BDE2B",
    9 => x"0023E92B",
    10 => x"007A64AE",
    11 => x"005FF480",
    12 => x"002F9A75",
    13 => x"0053DB0A",
    14 => x"002F7A49",
    15 => x"0028E527",
    16 => x"00299658",
    17 => x"000FA070",
    18 => x"006F65A5",
    19 => x"0036B788",
    20 => x"00777D91",
    21 => x"006ECAA1",
    22 => x"0027F968",
    23 => x"005FB37C",
    24 => x"005F8DD7",
    25 => x"0044FAE8",
    26 => x"006A84F8",
    27 => x"004DDC99",
    28 => x"001AD035",
    29 => x"007F9423",
    30 => x"003D3201",
    31 => x"000445C5",
    32 => x"00294A67",
    33 => x"00017620",
    34 => x"002EF4CD",
    35 => x"0035DEC5",
    36 => x"00668504",
    37 => x"0049102D",
    38 => x"005927D5",
    39 => x"003BBEAF",
    40 => x"0044F586",
    41 => x"00516E7D",
    42 => x"00368A96",
    43 => x"00541E42",
    44 => x"00360400",
    45 => x"007B4A4E",
    46 => x"0023D69C",
    47 => x"0077A55E",
    48 => x"0065F23E",
    49 => x"0066CAD7",
    50 => x"00357E1E",
    51 => x"00458F5A",
    52 => x"0035843F",
    53 => x"005F3618",
    54 => x"0067745D",
    55 => x"0038738C",
    56 => x"000C63A8",
    57 => x"00081B9A",
    58 => x"000E8F76",
    59 => x"003B3853",
    60 => x"003B8534",
    61 => x"0058DC31",
    62 => x"001F9D54",
    63 => x"00552F2E",
    64 => x"0043E6E6",
    65 => x"00688C82",
    66 => x"0047C1D0",
    67 => x"0051781A",
    68 => x"0069B65E",
    69 => x"003509EE",
    70 => x"002135C7",
    71 => x"0067AFBC",
    72 => x"006CAF76",
    73 => x"001D9772",
    74 => x"00419073",
    75 => x"00709CF7",
    76 => x"004F3281",
    77 => x"004FB2AF",
    78 => x"004870E1",
    79 => x"0001EFCA",
    80 => x"003410F2",
    81 => x"0070DE86",
    82 => x"0020C638",
    83 => x"00296E9F",
    84 => x"005297A4",
    85 => x"0047844C",
    86 => x"00799A6E",
    87 => x"005A140A",
    88 => x"0075A283",
    89 => x"006D2114",
    90 => x"007F863C",
    91 => x"006BE9F8",
    92 => x"007A0BDE",
    93 => x"001495D4",
    94 => x"001C4563",
    95 => x"006A0C63",
    96 => x"004CDBEA",
    97 => x"00040AF0",
    98 => x"0007C417",
    99 => x"002F4588",
    100 => x"0000AD00",
    101 => x"006F16BF",
    102 => x"000DCD44",
    103 => x"003C675A",
    104 => x"00470BCB",
    105 => x"007FBE7F",
    106 => x"00193948",
    107 => x"004E49C1",
    108 => x"0024756C",
    109 => x"007CA7E0",
    110 => x"000B98A1",
    111 => x"006BC809",
    112 => x"0002E46C",
    113 => x"0049A809",
    114 => x"003036C2",
    115 => x"00639FF7",
    116 => x"005B1C94",
    117 => x"007D2AE1",
    118 => x"00141305",
    119 => x"00147792",
    120 => x"00139E25",
    121 => x"0067B0E1",
    122 => x"00737945",
    123 => x"0069E803",
    124 => x"0051CEA3",
    125 => x"0044A79D",
    126 => x"00488058",
    127 => x"003A97D9",
    128 => x"001FEA93",
    129 => x"0033FF5A",
    130 => x"002358D4",
    131 => x"003A41F8",
    132 => x"004CDF73",
    133 => x"00223DFB",
    134 => x"005A8BA0",
    135 => x"00498423",
    136 => x"000412F5",
    137 => x"00252587",
    138 => x"006D04F1",
    139 => x"00359B5D",
    140 => x"004A28A1",
    141 => x"004682FD",
    142 => x"006D9B57",
    143 => x"004F25DF",
    144 => x"000DBE5E",
    145 => x"001C5E1A",
    146 => x"000DE0E6",
    147 => x"000C7F5A",
    148 => x"00078F83",
    149 => x"0067428B",
    150 => x"007F3705",
    151 => x"0077E6FD",
    152 => x"0075E022",
    153 => x"00503AF7",
    154 => x"001F0084",
    155 => x"0030EF86",
    156 => x"0049997E",
    157 => x"0077DCD7",
    158 => x"00742593",
    159 => x"004901C3",
    160 => x"00053919",
    161 => x"0004610C",
    162 => x"005AAD42",
    163 => x"003EB01B",
    164 => x"003472E7",
    165 => x"004CE03C",
    166 => x"001A7CC7",
    167 => x"00031924",
    168 => x"002B5EE5",
    169 => x"00291199",
    170 => x"00585A3B",
    171 => x"00134D71",
    172 => x"003DE11C",
    173 => x"00130984",
    174 => x"0025F051",
    175 => x"00185A46",
    176 => x"00466519",
    177 => x"001314BE",
    178 => x"00283891",
    179 => x"0049BB91",
    180 => x"0052308A",
    181 => x"001C853F",
    182 => x"001D0B4B",
    183 => x"006FD6A7",
    184 => x"006B88BF",
    185 => x"0012E11B",
    186 => x"004D3E3F",
    187 => x"006A0D30",
    188 => x"0078FDE5",
    189 => x"001406C7",
    190 => x"00327283",
    191 => x"0061ED6F",
    192 => x"006C5954",
    193 => x"001D4099",
    194 => x"00590579",
    195 => x"006AE5AE",
    196 => x"0016E405",
    197 => x"000BDBE7",
    198 => x"00221DE8",
    199 => x"0033F8CF",
    200 => x"00779935",
    201 => x"0054AA0D",
    202 => x"00665FF9",
    203 => x"0063B158",
    204 => x"0058711C",
    205 => x"00470C13",
    206 => x"000910D8",
    207 => x"00463E20",
    208 => x"00612659",
    209 => x"00251D8B",
    210 => x"002573B7",
    211 => x"007D5C90",
    212 => x"001DDD98",
    213 => x"00336898",
    214 => x"0002D4BB",
    215 => x"006D73A8",
    216 => x"004F4CBF",
    217 => x"00027C1C",
    218 => x"0018AA08",
    219 => x"002DFD71",
    220 => x"000C5CA5",
    221 => x"0019379A",
    222 => x"00478168",
    223 => x"00646C3E",
    224 => x"0051813D",
    225 => x"0035C539",
    226 => x"003B0115",
    227 => x"00041DC0",
    228 => x"0021C4F7",
    229 => x"0070FBF5",
    230 => x"001A35E7",
    231 => x"0007340E",
    232 => x"00795D46",
    233 => x"001A4CD0",
    234 => x"00645CAF",
    235 => x"001D2668",
    236 => x"00666E99",
    237 => x"006F0634",
    238 => x"007BE5DB",
    239 => x"00455FDC",
    240 => x"00530765",
    241 => x"005DC1B0",
    242 => x"007973DE",
    243 => x"005CFD0A",
    244 => x"0002CC93",
    245 => x"0070F806",
    246 => x"00189C2A",
    247 => x"0049C5AA",
    248 => x"00776A51",
    249 => x"003BCF2C",
    250 => x"007F234F",
    251 => x"006B16E0",
    252 => x"003C15CA",
    253 => x"00155E68",
    254 => x"0072F6B7",
    255 => x"001E29CE"
  );

begin
  sequential : process(clk)
  begin
    if (rising_edge(clk)) then
      --Read Logic
      q <= ram(to_integer(unsigned(address)));

    end if;
  end process;

end RTL;
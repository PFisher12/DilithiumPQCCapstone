library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use IEEE.math_real.all;
use work.GlobalVars.all;

entity bramTwoPort is
  generic (
    width   : integer := 32;
    depth   : integer := 8
  );

  	PORT
	(
    clk		      : IN STD_LOGIC;
		address_a		: IN STD_LOGIC_VECTOR (depth - 1 DOWNTO 0);
		address_b		: IN STD_LOGIC_VECTOR (depth - 1 DOWNTO 0);
		data_a		  : IN STD_LOGIC_VECTOR (width - 1 DOWNTO 0);
		data_b		  : IN STD_LOGIC_VECTOR (width - 1 DOWNTO 0);
		wren_a		  : IN STD_LOGIC  := '0';
		wren_b		  : IN STD_LOGIC  := '0';
		q_a		      : OUT STD_LOGIC_VECTOR (width - 1 DOWNTO 0);
		q_b		      : OUT STD_LOGIC_VECTOR (width - 1 DOWNTO 0)
	);

  attribute RAM_STYLE         : string;
  attribute RAM_STYLE of bramTwoPort : entity is "block";
end entity;

architecture RTL of bramTwoPort is
  subtype word_t is std_logic_vector(width - 1 downto 0);
  type memory_t is array(0 to 2**depth-1) of word_t;

  --shared variable ram : memory_t := (others => (others => '0'));
  shared variable ram : memory_t := (
    0 => x"006AAF4A",
    1 => x"000BC8BA",
    2 => x"004A1708",
    3 => x"0069EF16",
    4 => x"000E9F72",
    5 => x"00750878",
    6 => x"00628125",
    7 => x"0063AF19",
    8 => x"000EDD20",
    9 => x"005074A2",
    10 => x"006AF77B",
    11 => x"0022F600",
    12 => x"00416CB5",
    13 => x"005535DC",
    14 => x"005093DB",
    15 => x"00586CBE",
    16 => x"003420E5",
    17 => x"0058368F",
    18 => x"000D3705",
    19 => x"00093A4C",
    20 => x"006B3F95",
    21 => x"0046F780",
    22 => x"007B4E4D",
    23 => x"0025B5C1",
    24 => x"00422E40",
    25 => x"0002CDF9",
    26 => x"002D2E1A",
    27 => x"00600925",
    28 => x"00260262",
    29 => x"002F2310",
    30 => x"0022310F",
    31 => x"0053EF51",
    32 => x"007073D7",
    33 => x"00565F03",
    34 => x"0020CEA2",
    35 => x"00785931",
    36 => x"005F3643",
    37 => x"007511AA",
    38 => x"0038E982",
    39 => x"00639102",
    40 => x"006751FB",
    41 => x"006304C9",
    42 => x"003B9016",
    43 => x"0035EBAC",
    44 => x"000F7241",
    45 => x"00410C84",
    46 => x"0020F078",
    47 => x"0031D1D4",
    48 => x"001D3369",
    49 => x"005E49B2",
    50 => x"0028080B",
    51 => x"0045198F",
    52 => x"004601BD",
    53 => x"003DAC22",
    54 => x"005ECA2E",
    55 => x"001FF952",
    56 => x"0006718C",
    57 => x"001CD4E1",
    58 => x"004E50D6",
    59 => x"004061F3",
    60 => x"007C4302",
    61 => x"00116D9D",
    62 => x"0006B5B5",
    63 => x"00752648",
    64 => x"0009C3C5",
    65 => x"001DA3EF",
    66 => x"0058D930",
    67 => x"00588603",
    68 => x"001C7AE8",
    69 => x"000086EE",
    70 => x"00755591",
    71 => x"00124E60",
    72 => x"004E2527",
    73 => x"000B4098",
    74 => x"0075BEF0",
    75 => x"0024EBEB",
    76 => x"0043DD9E",
    77 => x"005FBD1A",
    78 => x"0060F998",
    79 => x"005C7B4E",
    80 => x"00283FC8",
    81 => x"0071810C",
    82 => x"00609DF5",
    83 => x"00714814",
    84 => x"0016337B",
    85 => x"007267FB",
    86 => x"0015716F",
    87 => x"0062A3C6",
    88 => x"004D68D6",
    89 => x"00620792",
    90 => x"000EDCA4",
    91 => x"001EAEAC",
    92 => x"003961A1",
    93 => x"00316F4C",
    94 => x"0038A224",
    95 => x"002F88EA",
    96 => x"0001E3CA",
    97 => x"0030539D",
    98 => x"005311C6",
    99 => x"0079814E",
    100 => x"005B2F16",
    101 => x"003454DB",
    102 => x"0077A3A5",
    103 => x"000C6335",
    104 => x"007A479F",
    105 => x"003DF54B",
    106 => x"0016406D",
    107 => x"003F2A0A",
    108 => x"007825A5",
    109 => x"004917CD",
    110 => x"00285AAF",
    111 => x"001B525C",
    112 => x"002FBD9C",
    113 => x"002492B4",
    114 => x"00518AD2",
    115 => x"005E68E3",
    116 => x"0029377B",
    117 => x"0027C78E",
    118 => x"007ED20F",
    119 => x"0042406C",
    120 => x"006C7EDD",
    121 => x"00485761",
    122 => x"004E19ED",
    123 => x"00118534",
    124 => x"005F97F8",
    125 => x"002EFBA9",
    126 => x"00153606",
    127 => x"007CF316",
    128 => x"0032A53D",
    129 => x"006C2E23",
    130 => x"00362EB0",
    131 => x"003481D3",
    132 => x"007B4F1C",
    133 => x"004D6054",
    134 => x"0012AE45",
    135 => x"004603D8",
    136 => x"00712F1B",
    137 => x"005F2EDC",
    138 => x"004562DB",
    139 => x"002B251E",
    140 => x"00002D22",
    141 => x"0030EED5",
    142 => x"004ECA1F",
    143 => x"001694CE",
    144 => x"007AFCA7",
    145 => x"004AFC19",
    146 => x"0048B3C6",
    147 => x"002642DD",
    148 => x"00440420",
    149 => x"0026AD33",
    150 => x"007D7D07",
    151 => x"0050D1D4",
    152 => x"001BB903",
    153 => x"004650F3",
    154 => x"001E7EC0",
    155 => x"005DC155",
    156 => x"0035BB1A",
    157 => x"000A31EC",
    158 => x"0045DB55",
    159 => x"0025E1EC",
    160 => x"000635AD",
    161 => x"007A0FB3",
    162 => x"005F5319",
    163 => x"007DD5E4",
    164 => x"0027824E",
    165 => x"003ED4A9",
    166 => x"00165063",
    167 => x"0067DB5F",
    168 => x"001CBEE3",
    169 => x"006361E9",
    170 => x"00206EE2",
    171 => x"0041A9FC",
    172 => x"003884B5",
    173 => x"00274858",
    174 => x"004E15F6",
    175 => x"003FBD95",
    176 => x"002FC8D2",
    177 => x"0027B20E",
    178 => x"002DB714",
    179 => x"0077B129",
    180 => x"007A0DB9",
    181 => x"00431A03",
    182 => x"0023F99C",
    183 => x"001B4EE0",
    184 => x"003BC38C",
    185 => x"000241AD",
    186 => x"007B7A90",
    187 => x"0057151A",
    188 => x"0011594E",
    189 => x"002B47A4",
    190 => x"001B3359",
    191 => x"0035321B",
    192 => x"00032E71",
    193 => x"006F2779",
    194 => x"0022EEE8",
    195 => x"007535D9",
    196 => x"0008C89A",
    197 => x"00105325",
    198 => x"00488C4A",
    199 => x"000986D5",
    200 => x"00538D2F",
    201 => x"007C2FBC",
    202 => x"004B8C6F",
    203 => x"00339870",
    204 => x"001D1207",
    205 => x"002B9BDB",
    206 => x"002473D3",
    207 => x"0047EDBD",
    208 => x"006129C1",
    209 => x"0053B7AF",
    210 => x"0052565F",
    211 => x"0013272B",
    212 => x"006CEBBA",
    213 => x"003181EE",
    214 => x"003657B5",
    215 => x"000C581F",
    216 => x"005F1EE8",
    217 => x"0019B205",
    218 => x"0051510E",
    219 => x"00724791",
    220 => x"007B569F",
    221 => x"0036886F",
    222 => x"007C7AD7",
    223 => x"000CB5EC",
    224 => x"0046802F",
    225 => x"003E9712",
    226 => x"0019224F",
    227 => x"003A6264",
    228 => x"002C370C",
    229 => x"00100F2A",
    230 => x"00574C25",
    231 => x"006B5FED",
    232 => x"0060BD5D",
    233 => x"0079C32E",
    234 => x"004460A0",
    235 => x"000A37D0",
    236 => x"00499DCB",
    237 => x"00126EB8",
    238 => x"003BF4BB",
    239 => x"00081D82",
    240 => x"006883B2",
    241 => x"006D5B70",
    242 => x"006F300F",
    243 => x"005C79C9",
    244 => x"002AE1BA",
    245 => x"000F9971",
    246 => x"0048300F",
    247 => x"001B3E51",
    248 => x"00138999",
    249 => x"00770790",
    250 => x"0028B38D",
    251 => x"001335BD",
    252 => x"0052CD98",
    253 => x"007F95AE",
    254 => x"0046E9FB",
    255 => x"006419C6");


begin

  

  sequential1 : process(clk)
  begin
    if (clk'event and clk = '1') then
      --Write Logic
      if(wren_a = '1') then
        ram(to_integer(unsigned(address_a))) := data_a;
      end if;
      --Read Logic
      q_a <= ram(to_integer(unsigned(address_a)));
    end if;
  end process;


  sequential2 : process(clk)
  begin
    if (clk'event and clk = '1') then
      --Write Logic
      if(wren_b = '1') then
        ram(to_integer(unsigned(address_b))) := data_b;
      end if;
      --Read Logic
      q_b <= ram(to_integer(unsigned(address_b)));
    end if;
  end process;


end RTL;
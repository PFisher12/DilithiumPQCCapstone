library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use IEEE.math_real.all;
use work.GlobalVars.all;

entity romInverseZetas is
  generic (
    width   : integer := 32;
    depth   : integer := 8
  );

  	PORT
	(
		address 		: IN STD_LOGIC_VECTOR (depth - 1 DOWNTO 0);
		clk		    : IN STD_LOGIC;
		q		        : OUT STD_LOGIC_VECTOR (width - 1 DOWNTO 0)
	);

  attribute RAM_STYLE         : string;
  attribute RAM_STYLE of romInverseZetas : entity is "block";
end entity;

architecture RTL of romInverseZetas is
  subtype word_t is std_logic_vector(width - 1 downto 0);
  type memory_t is array(0 to 2**depth-1) of word_t;

  signal ram : memory_t := (
    0 => x"0061B633",
    1 => x"000CE94A",
    2 => x"006A8199",
    3 => x"0043CA37",
    4 => x"0014C921",
    5 => x"0000BCB2",
    6 => x"004410D5",
    7 => x"000875B0",
    8 => x"00361A57",
    9 => x"006743D7",
    10 => x"000EE7FB",
    11 => x"007D136E",
    12 => x"0022E2F7",
    13 => x"00066C23",
    14 => x"00221E51",
    15 => x"002CD89C",
    16 => x"003A8025",
    17 => x"0003FA26",
    18 => x"0010D9CD",
    19 => x"00197168",
    20 => x"0062B999",
    21 => x"001B8352",
    22 => x"00659331",
    23 => x"000682BB",
    24 => x"0078ABF3",
    25 => x"0065AA1A",
    26 => x"000EE40C",
    27 => x"005E1B0A",
    28 => x"007BC241",
    29 => x"0044DEEC",
    30 => x"004A1AC8",
    31 => x"002E5EC4",
    32 => x"001B73C3",
    33 => x"00385E99",
    34 => x"0066A867",
    35 => x"0073835C",
    36 => x"0051E290",
    37 => x"006735F9",
    38 => x"007D63E5",
    39 => x"00309342",
    40 => x"00126C59",
    41 => x"007D0B46",
    42 => x"004C7769",
    43 => x"00620269",
    44 => x"00028371",
    45 => x"005A6C4A",
    46 => x"005AC276",
    47 => x"001EB9A8",
    48 => x"0039A1E1",
    49 => x"0076CF29",
    50 => x"0038D3EE",
    51 => x"00276EE5",
    52 => x"001C2EA9",
    53 => x"00198008",
    54 => x"002B35F4",
    55 => x"000846CC",
    56 => x"004BE732",
    57 => x"005DC219",
    58 => x"0074041A",
    59 => x"0068FBFC",
    60 => x"0014FA53",
    61 => x"0026DA88",
    62 => x"00629F68",
    63 => x"001386AD",
    64 => x"001DF292",
    65 => x"004D6D7E",
    66 => x"006BD93A",
    67 => x"0006E21C",
    68 => x"0015D2D1",
    69 => x"0032A1C2",
    70 => x"006CFEE6",
    71 => x"00145742",
    72 => x"0010095A",
    73 => x"0062D4B6",
    74 => x"00635AC2",
    75 => x"002DAF77",
    76 => x"00362470",
    77 => x"0057A770",
    78 => x"006CCB43",
    79 => x"00397AE8",
    80 => x"006785BB",
    81 => x"0059EFB0",
    82 => x"006CD67D",
    83 => x"0041FEE5",
    84 => x"006C9290",
    85 => x"002785C6",
    86 => x"0056CE68",
    87 => x"0054811C",
    88 => x"007CC6DD",
    89 => x"0065633A",
    90 => x"0032FFC5",
    91 => x"004B6D1A",
    92 => x"00412FE6",
    93 => x"002532BF",
    94 => x"007B7EF5",
    95 => x"007AA6E8",
    96 => x"0036DE3E",
    97 => x"000BBA6E",
    98 => x"0008032A",
    99 => x"00364683",
    100 => x"004EF07B",
    101 => x"0060DF7D",
    102 => x"002FA50A",
    103 => x"0009FFDF",
    104 => x"0007F904",
    105 => x"0000A8FC",
    106 => x"00189D76",
    107 => x"0078507E",
    108 => x"007360A7",
    109 => x"0071FF1B",
    110 => x"006381E7",
    111 => x"007221A3",
    112 => x"0030BA22",
    113 => x"001244AA",
    114 => x"00395D04",
    115 => x"0035B760",
    116 => x"004A44A4",
    117 => x"0012DB10",
    118 => x"005ABA7A",
    119 => x"007BCD0C",
    120 => x"00365BDE",
    121 => x"00255461",
    122 => x"005DA206",
    123 => x"0033008E",
    124 => x"00459E09",
    125 => x"005C872D",
    126 => x"004BE0A7",
    127 => x"005FF56E",
    128 => x"00454828",
    129 => x"00375FA9",
    130 => x"003B3864",
    131 => x"002E115E",
    132 => x"0015F7FE",
    133 => x"000C66BC",
    134 => x"00182F20",
    135 => x"006C41DC",
    136 => x"006B686F",
    137 => x"006BCCFC",
    138 => x"0002B520",
    139 => x"0024C36D",
    140 => x"001C400A",
    141 => x"004FA93F",
    142 => x"003637F8",
    143 => x"007CFB95",
    144 => x"001417F8",
    145 => x"00744760",
    146 => x"00033821",
    147 => x"005B6A95",
    148 => x"00319640",
    149 => x"0066A6B9",
    150 => x"00002182",
    151 => x"0038D436",
    152 => x"004378A7",
    153 => x"007212BD",
    154 => x"0010C942",
    155 => x"007F3301",
    156 => x"00509A79",
    157 => x"00781BEA",
    158 => x"007BD511",
    159 => x"00330417",
    160 => x"0015D39E",
    161 => x"00639A9E",
    162 => x"006B4A2D",
    163 => x"0005D423",
    164 => x"0013F609",
    165 => x"000059C5",
    166 => x"0012BEED",
    167 => x"000A3D7E",
    168 => x"0025CBF7",
    169 => x"00064593",
    170 => x"00385BB5",
    171 => x"002D485D",
    172 => x"00567162",
    173 => x"005F19C9",
    174 => x"000F017B",
    175 => x"004BCF0F",
    176 => x"007DF037",
    177 => x"00376F20",
    178 => x"00302D52",
    179 => x"0030AD80",
    180 => x"000F430A",
    181 => x"003E4F8E",
    182 => x"0062488F",
    183 => x"0013308B",
    184 => x"00183045",
    185 => x"005EAA3A",
    186 => x"004AD613",
    187 => x"001629A3",
    188 => x"002E67E7",
    189 => x"00381E31",
    190 => x"0017537F",
    191 => x"003BF91B",
    192 => x"002AB0D3",
    193 => x"006042AD",
    194 => x"002703D0",
    195 => x"00445ACD",
    196 => x"0044A7AE",
    197 => x"0071508B",
    198 => x"0077C467",
    199 => x"00737C59",
    200 => x"00476C75",
    201 => x"00186BA4",
    202 => x"0020A9E9",
    203 => x"004A5BC2",
    204 => x"003A50A7",
    205 => x"004A61E3",
    206 => x"0019152A",
    207 => x"0019EDC3",
    208 => x"00083AA3",
    209 => x"005C0965",
    210 => x"000495B3",
    211 => x"0049DC01",
    212 => x"002BC1BF",
    213 => x"0049556B",
    214 => x"002E7184",
    215 => x"003AEA7B",
    216 => x"00442152",
    217 => x"0026B82C",
    218 => x"0036CFD4",
    219 => x"00195AFD",
    220 => x"004A013C",
    221 => x"0050EB34",
    222 => x"007E69E1",
    223 => x"0056959A",
    224 => x"007B9A3C",
    225 => x"0042AE00",
    226 => x"00004BDE",
    227 => x"00650FCC",
    228 => x"00320368",
    229 => x"00155B09",
    230 => x"003AE519",
    231 => x"0020522A",
    232 => x"00202C85",
    233 => x"0057E699",
    234 => x"00111560",
    235 => x"00086270",
    236 => x"00492879",
    237 => x"00107A5C",
    238 => x"00703F91",
    239 => x"005649A9",
    240 => x"0056FADA",
    241 => x"005065B8",
    242 => x"002C04F7",
    243 => x"0050458C",
    244 => x"001FEB81",
    245 => x"00057B53",
    246 => x"005BF6D6",
    247 => x"006401D6",
    248 => x"0078C1DD",
    249 => x"000D5ED8",
    250 => x"000BDEE8",
    251 => x"007C41BD",
    252 => x"0007EAFD",
    253 => x"0027CEFE",
    254 => x"007F7B0A",
    255 => x"00000000"
  );

begin
  sequential : process(clk)
  begin
    if (rising_edge(clk)) then
      --Read Logic
      q <= ram(to_integer(unsigned(address)));

    end if;
  end process;

end RTL;